module qoi
