module qoi

